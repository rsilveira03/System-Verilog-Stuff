module top;
	int a = 10;
	initial begin
		$display(a = %0d",a);
	end
endmodule